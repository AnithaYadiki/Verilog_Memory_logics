module clk_buff(input mclk,output bclk);

buf buff(bclk,mclk);

endmodule
